grammar edu:umn:cs:melt:dcv2:monto;
